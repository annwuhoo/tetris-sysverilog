//Sprite Table for Expansion by Factor
//Single block is a 4x4 block for Acting Blocks
//Single block in TETRIS font is 8x8 block
//These factors can be changed in the ColorMapper under varaibles fe and te respectively
module Sprite_Table_FE (
					// variable [#Cols][#Rows][EntryDepth]
					 output logic [4:0][22:0][3:0] HOLD,
					 output logic [4:0][30:0][3:0] ANNWU,
					 output logic [4:0][53:0][3:0] PATRICKSU,
					 output logic [10:0][24:0][3:0] GAMEOVER,
					 output logic [4:0][39:0][3:0] TETRIS_h,
					 output logic [39:0][4:0][3:0] TETRIS,
					 output logic [39:0][4:0][3:0] TETRIS2,
					 output logic [3:0][15:0][3:0] I_block_h,
					 output logic [15:0][3:0][3:0] I_block_v,
					 output logic [7:0][7:0][3:0] O_block,
					 output logic [7:0][11:0][3:0] J_block_0,
					 output logic [11:0][7:0][3:0] J_block_1,
					 output logic [7:0][11:0][3:0] J_block_2,
					 output logic [11:0][7:0][3:0] J_block_3,
					 output logic [7:0][11:0][3:0] T_block_0,
					 output logic [11:0][7:0][3:0] T_block_1,
					 output logic [7:0][11:0][3:0] T_block_2,
					 output logic [11:0][7:0][3:0] T_block_3,
					 output logic [7:0][11:0][3:0] L_block_0,
					 output logic [11:0][7:0][3:0] L_block_1,
					 output logic [7:0][11:0][3:0] L_block_2,
					 output logic [11:0][7:0][3:0] L_block_3,
					 output logic [7:0][11:0][3:0] S_block_0,
					 output logic [11:0][7:0][3:0] S_block_1,
					 output logic [7:0][11:0][3:0] Z_block_0,
					 output logic [11:0][7:0][3:0] Z_block_1,
					 output logic [4:0][28:0][3:0] SCORE_Letters,
					 output logic [4:0][4:0][3:0] zero,
					 output logic [4:0][4:0][3:0] one,
					 output logic [4:0][4:0][3:0] two,
					 output logic [4:0][4:0][3:0] three,
					 output logic [4:0][4:0][3:0] four,
					 output logic [4:0][4:0][3:0] five,
					 output logic [4:0][4:0][3:0] six,
					 output logic [4:0][4:0][3:0] seven,
					 output logic [4:0][4:0][3:0] eight,
					 output logic [4:0][4:0][3:0] nine);
	 
	//Single Standard Block is 16x16
	always_comb
	begin
	
	I_block_h <= '{
	
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,1,1,7,7,1,1,7,7,1,1,7,7,1,1,7},
		'{7,1,1,7,7,1,1,7,7,1,1,7,7,1,1,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}
	};
	
	I_block_v <= '{
		
		'{7,7,7,7},
		'{7,1,1,7},
		'{7,1,1,7},
		'{7,7,7,7},
		'{7,7,7,7},
		'{7,1,1,7},
		'{7,1,1,7},
		'{7,7,7,7},
		'{7,7,7,7},
		'{7,1,1,7},
		'{7,1,1,7},
		'{7,7,7,7},
		'{7,7,7,7},
		'{7,1,1,7},
		'{7,1,1,7},
		'{7,7,7,7}
	};


	O_block <= '{
	
		'{7,7,7,7,7,7,7,7},
		'{7,2,2,7,7,2,2,7},
		'{7,2,2,7,7,2,2,7},
		'{7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7},
		'{7,2,2,7,7,2,2,7},
		'{7,2,2,7,7,2,2,7},
		'{7,7,7,7,7,7,7,7}
	};
	
	J_block_0 <= '{
	
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,3,3,7,7,3,3,7,7,3,3,7},
		'{7,3,3,7,7,3,3,7,7,3,3,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7},
		'{0,0,0,0,0,0,0,0,7,7,7,7},
		'{0,0,0,0,0,0,0,0,7,3,3,7},
		'{0,0,0,0,0,0,0,0,7,3,3,7},
		'{0,0,0,0,0,0,0,0,7,7,7,7}
	};
	
	J_block_1 <= '{
	
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,3,3,7},
	'{0,0,0,0,7,3,3,7},
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,3,3,7},
	'{0,0,0,0,7,3,3,7},
	'{0,0,0,0,7,7,7,7},
	'{7,7,7,7,7,7,7,7},
	'{7,3,3,7,7,3,3,7},
	'{7,3,3,7,7,3,3,7},
	'{7,7,7,7,7,7,7,7}
	};
	
	J_block_2 <= '{
	
	'{7,7,7,7,0,0,0,0,0,0,0,0},
	'{7,3,3,7,0,0,0,0,0,0,0,0},
	'{7,3,3,7,0,0,0,0,0,0,0,0},
	'{7,7,7,7,0,0,0,0,0,0,0,0},
	'{7,7,7,7,7,7,7,7,7,7,7,7},
	'{7,3,3,7,7,3,3,7,7,3,3,7},
	'{7,3,3,7,7,3,3,7,7,3,3,7},
	'{7,7,7,7,7,7,7,7,7,7,7,7}
	};

	J_block_3 <= '{
	
	'{7,7,7,7,7,7,7,7},
	'{7,3,3,7,7,3,3,7},
	'{7,3,3,7,7,3,3,7},
	'{7,7,7,7,7,7,7,7},
	'{7,7,7,7,0,0,0,0},
	'{7,3,3,7,0,0,0,0},
	'{7,3,3,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0},
	'{7,3,3,7,0,0,0,0},
	'{7,3,3,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0}
	};
	
	L_block_0 <= ' {
	
	'{7,7,7,7,7,7,7,7,7,7,7,7},
	'{7,4,4,7,7,4,4,7,7,4,4,7},
	'{7,4,4,7,7,4,4,7,7,4,4,7},
	'{7,7,7,7,7,7,7,7,7,7,7,7},
	'{7,7,7,7,0,0,0,0,0,0,0,0},
	'{7,4,4,7,0,0,0,0,0,0,0,0},
	'{7,4,4,7,0,0,0,0,0,0,0,0},
	'{7,7,7,7,0,0,0,0,0,0,0,0}
	
	};

	L_block_1 <= ' {
	
	'{7,7,7,7,7,7,7,7},
	'{7,4,4,7,7,4,4,7},
	'{7,4,4,7,7,4,4,7},
	'{7,7,7,7,7,7,7,7},
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,4,4,7},
	'{0,0,0,0,7,4,4,7},
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,4,4,7},
	'{0,0,0,0,7,4,4,7},
	'{0,0,0,0,7,7,7,7}
	};

	L_block_2 <= ' {
	
  '{0,0,0,0,0,0,0,0,7,7,7,7},
  '{0,0,0,0,0,0,0,0,7,4,4,7},
  '{0,0,0,0,0,0,0,0,7,4,4,7},
  '{0,0,0,0,0,0,0,0,7,7,7,7},
  '{7,7,7,7,7,7,7,7,7,7,7,7},
  '{7,4,4,7,7,4,4,7,7,4,4,7},
  '{7,4,4,7,7,4,4,7,7,4,4,7},
  '{7,7,7,7,7,7,7,7,7,7,7,7}
	
	};

	L_block_3 <= ' {
	
	'{7,7,7,7,0,0,0,0},
	'{7,4,4,7,0,0,0,0},
	'{7,4,4,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0},
	'{7,4,4,7,0,0,0,0},
	'{7,4,4,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0},
	'{7,7,7,7,7,7,7,7},
	'{7,4,4,7,7,4,4,7},
	'{7,4,4,7,7,4,4,7},
	'{7,7,7,7,7,7,7,7}	
	};
	
	S_block_0 <= '{
	
	'{0,0,0,0,7,7,7,7,7,7,7,7},
	'{0,0,0,0,7,5,5,7,7,5,5,7},
	'{0,0,0,0,7,5,5,7,7,5,5,7},
	'{0,0,0,0,7,7,7,7,7,7,7,7},
	'{7,7,7,7,7,7,7,7,0,0,0,0},
	'{7,5,5,7,7,5,5,7,0,0,0,0},
	'{7,5,5,7,7,5,5,7,0,0,0,0},
	'{7,7,7,7,7,7,7,7,0,0,0,0}
	};
	
	S_block_1 <= '{
	
	'{7,7,7,7,0,0,0,0},
	'{7,5,5,7,0,0,0,0},
	'{7,5,5,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0},
	'{7,7,7,7,7,7,7,7},
	'{7,5,5,7,7,5,5,7},
	'{7,5,5,7,7,5,5,7},
	'{7,7,7,7,7,7,7,7},
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,5,5,7},
	'{0,0,0,0,7,5,5,7},
	'{0,0,0,0,7,7,7,7}
	};
	
	Z_block_0 <= '{
	
	'{7,7,7,7,7,7,7,7,0,0,0,0},
	'{7,6,6,7,7,6,6,7,0,0,0,0},
	'{7,6,6,7,7,6,6,7,0,0,0,0},
	'{7,7,7,7,7,7,7,7,0,0,0,0},
	'{0,0,0,0,7,7,7,7,7,7,7,7},
	'{0,0,0,0,7,6,6,7,7,6,6,7},
	'{0,0,0,0,7,6,6,7,7,6,6,7},
	'{0,0,0,0,7,7,7,7,7,7,7,7}	
	
	};
	
	Z_block_1 <= '{
	
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,6,6,7},
	'{0,0,0,0,7,6,6,7},
	'{0,0,0,0,7,7,7,7},
	'{7,7,7,7,7,7,7,7},
	'{7,6,6,7,7,6,6,7},
	'{7,6,6,7,7,6,6,7},
	'{7,7,7,7,7,7,7,7},
	'{7,7,7,7,0,0,0,0},
	'{7,6,6,7,0,0,0,0},
	'{7,6,6,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0}
	
	};
	
	T_block_0 <= '{
	
	'{7,7,7,7,7,7,7,7,7,7,7,7},
	'{7,8,8,7,7,8,8,7,7,8,8,7},
	'{7,8,8,7,7,8,8,7,7,8,8,7},
	'{7,7,7,7,7,7,7,7,7,7,7,7},
	'{0,0,0,0,7,7,7,7,0,0,0,0},
	'{0,0,0,0,7,8,8,7,0,0,0,0},
	'{0,0,0,0,7,8,8,7,0,0,0,0},
	'{0,0,0,0,7,7,7,7,0,0,0,0}
	
	};
	
	T_block_1 <= '{
	
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,8,8,7},
	'{0,0,0,0,7,8,8,7},
	'{0,0,0,0,7,7,7,7},
	'{7,7,7,7,7,7,7,7},
	'{7,8,8,7,7,8,8,7},
	'{7,8,8,7,7,8,8,7},
	'{7,7,7,7,7,7,7,7},
	'{0,0,0,0,7,7,7,7},
	'{0,0,0,0,7,8,8,7},
	'{0,0,0,0,7,8,8,7},
	'{0,0,0,0,7,7,7,7}
	
	};
	
	T_block_2 <= '{
	
	'{0,0,0,0,7,7,7,7,0,0,0,0},
	'{0,0,0,0,7,8,8,7,0,0,0,0},
	'{0,0,0,0,7,8,8,7,0,0,0,0},
	'{0,0,0,0,7,7,7,7,0,0,0,0},
	'{7,7,7,7,7,7,7,7,7,7,7,7},
	'{7,8,8,7,7,8,8,7,7,8,8,7},
	'{7,8,8,7,7,8,8,7,7,8,8,7},
	'{7,7,7,7,7,7,7,7,7,7,7,7}
	
	};
	
	T_block_3 <= '{
	
	'{7,7,7,7,0,0,0,0},
	'{7,8,8,7,0,0,0,0},
	'{7,8,8,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0},
	'{7,7,7,7,7,7,7,7},
	'{7,8,8,7,7,8,8,7},
	'{7,8,8,7,7,8,8,7},
	'{7,7,7,7,7,7,7,7},
	'{7,7,7,7,0,0,0,0},
	'{7,8,8,7,0,0,0,0},
	'{7,8,8,7,0,0,0,0},
	'{7,7,7,7,0,0,0,0}
	
	};
//UPSIDE DOWN
TETRIS <= '{
	'{0,0,0,0,0},
	'{0,0,0,0,0},
	'{0,0,0,0,0},
	'{6,6,6,6,6},
	'{0,0,6,0,0},
	'{0,0,6,0,0},
	'{0,0,6,0,0},
	'{0,0,6,0,0},
	'{0,0,0,0,0},
	'{4,4,4,4,4},
	'{4,0,0,0,0},
	'{4,4,4,4,4},
	'{4,0,0,0,0},
	'{4,4,4,4,4},
	'{0,0,0,0,0},
	'{2,2,2,2,2},
	'{0,0,2,0,0},
	'{0,0,2,0,0},
	'{0,0,2,0,0},
	'{0,0,2,0,0},
	'{0,0,0,0,0},
	'{5,5,5,5,5},
	'{5,0,0,0,5},
	'{5,5,5,5,5},
	'{5,0,0,5,0},
	'{5,0,0,0,5},
	'{0,0,0,0,0},
	'{1,1,1,1,1},
	'{0,0,1,0,0},
	'{0,0,1,0,0},
	'{0,0,1,0,0},
	'{1,1,1,1,1},
	'{0,0,0,0,0},
	'{8,8,8,8,8},
	'{8,0,0,0,0},
	'{8,8,8,8,8},
	'{0,0,0,0,8},
	'{8,8,8,8,8},
	'{0,0,0,0,0},
	'{0,0,0,0,0}
};

//RIGHTSIDE UP
TETRIS2 <= '{
	'{0,0,0,0,0},
	'{0,0,0,0,0},
	'{0,0,0,0,0},
	'{8,8,8,8,8},
	'{8,0,0,0,0},
	'{8,8,8,8,8},
	'{0,0,0,0,8},
	'{8,8,8,8,8},
	'{0,0,0,0,0},
	'{1,1,1,1,1},
	'{0,0,1,0,0},
	'{0,0,1,0,0},
	'{0,0,1,0,0},
	'{1,1,1,1,1},
	'{0,0,0,0,0},
	'{5,0,0,0,5},
	'{0,5,0,0,5},
	'{5,5,5,5,5},
	'{5,0,0,0,5},
	'{5,5,5,5,5},
	'{0,0,0,0,0},
	'{0,0,2,0,0},
	'{0,0,2,0,0},
	'{0,0,2,0,0},
	'{0,0,2,0,0},
	'{2,2,2,2,2},
	'{0,0,0,0,0},
	'{4,4,4,4,4},
	'{0,0,0,0,4},
	'{4,4,4,4,4},
	'{0,0,0,0,4},
	'{4,4,4,4,4},
	'{0,0,0,0,0},
	'{0,0,6,0,0},
	'{0,0,6,0,0},
	'{0,0,6,0,0},
	'{0,0,6,0,0},
	'{6,6,6,6,6},
	'{0,0,0,0,0},
	'{0,0,0,0,0}
};

TETRIS_h <= '{
	
		'{0,0,8,8,8,8,8,0,1,1,1,1,1,0,5,0,0,0,5,0,0,0,2,0,0,0,4,4,4,4,4,0,0,0,6,0,0,0,0,0},
		'{0,0,8,0,0,0,0,0,0,0,1,0,0,0,0,5,0,0,5,0,0,0,2,0,0,0,0,0,0,0,4,0,0,0,6,0,0,0,0,0},
		'{0,0,8,8,8,8,8,0,0,0,1,0,0,0,5,5,5,5,5,0,0,0,2,0,0,0,4,4,4,4,4,0,0,0,6,0,0,0,0,0},
		'{0,0,0,0,0,0,8,0,0,0,1,0,0,0,5,0,0,0,5,0,0,0,2,0,0,0,0,0,0,0,4,0,0,0,6,0,0,0,0,0},
		'{0,0,8,8,8,8,8,0,1,1,1,1,1,0,5,5,5,5,5,0,2,2,2,2,2,0,4,4,4,4,4,0,6,6,6,6,6,0,0,0}
		
	};
	
	GAMEOVER <= '{
	
'{0,4,0,0,0,4,0,6,6,6,6,6,0,0,0,8,0,0,0,1,1,1,1,1,0},
'{0,0,4,0,0,4,0,0,0,0,0,6,0,8,8,0,8,8,0,1,0,0,0,1,0},
'{0,4,4,4,4,4,0,6,6,6,6,6,0,8,0,0,0,8,0,1,0,0,0,1,0},
'{0,4,0,0,0,4,0,0,0,0,0,6,0,8,0,0,0,8,0,1,0,0,0,1,0},
'{0,4,4,4,4,4,0,6,6,6,6,6,0,8,0,0,0,8,0,1,1,1,1,1,0},
'{0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
'{0,5,5,5,5,5,0,2,0,0,0,2,0,4,0,0,0,4,0,6,6,6,6,6,0},
'{0,0,0,0,0,5,0,2,0,0,0,2,0,4,0,0,0,4,0,6,0,0,0,6,0},
'{0,5,5,5,5,5,0,2,0,2,0,2,0,4,4,4,4,4,0,6,6,0,0,6,0},
'{0,0,0,0,0,5,0,2,2,0,2,2,0,4,0,0,0,4,0,0,0,0,0,6,0},
'{0,5,5,5,5,5,0,2,0,0,0,2,0,4,4,4,4,4,0,6,6,6,6,6,0}

};
	SCORE_Letters <= '{
	
	'{4,4,4,4,4,0,2,0,0,0,2,0,5,5,5,5,5,0,1,1,1,1,1,0,8,8,8,8,8},
	'{0,0,0,0,4,0,0,2,0,0,2,0,5,0,0,0,5,0,0,0,0,0,1,0,8,0,0,0,0},
	'{4,4,4,4,4,0,2,2,2,2,2,0,5,0,0,0,5,0,0,0,0,0,1,0,8,8,8,8,8},
	'{0,0,0,0,4,0,2,0,0,0,2,0,5,0,0,0,5,0,0,0,0,0,1,0,0,0,0,0,8},
	'{4,4,4,4,4,0,2,2,2,2,2,0,5,5,5,5,5,0,1,1,1,1,1,0,8,8,8,8,8}
	
	};
	
	
HOLD <= '{

 '{0,1,1,1,1,0,5,5,5,5,5,0,2,2,2,2,2,0,4,0,0,0,4},
 '{1,0,0,0,1,0,0,0,0,0,5,0,2,0,0,0,2,0,4,0,0,0,4},
 '{1,0,0,0,1,0,0,0,0,0,5,0,2,0,0,0,2,0,4,4,4,4,4},
 '{1,0,0,0,1,0,0,0,0,0,5,0,2,0,0,0,2,0,4,0,0,0,4},
 '{0,1,1,1,1,0,0,0,0,0,5,0,2,2,2,2,2,0,4,0,0,0,4}
 
 };


	zero <= '{
	
	'{9,9,9,9,9},
	'{9,0,0,0,9},
	'{9,0,0,0,9},
	'{9,0,0,0,9},
	'{9,9,9,9,9}

};
	
	
	one <= '{
	
	'{0,0,9,0,0},
	'{0,0,9,0,0},
	'{0,0,9,0,0},
	'{0,0,9,0,0},
	'{0,0,9,0,0}
	
	};	
	
	two <= '{

	'{9,9,9,9,9},
	'{0,0,0,0,9},
	'{9,9,9,9,9},
	'{9,0,0,0,0},
	'{9,9,9,9,9}
	
	};

	three <= '{
	
	'{9,9,9,9,9},
	'{9,0,0,0,0},
	'{9,9,9,9,9},
	'{9,0,0,0,0},
	'{9,9,9,9,9}
};
	
	
	
	four <= '{
	
	'{9,0,0,0,0},
	'{9,0,0,0,0},
	'{9,9,9,9,9},
	'{9,0,0,0,9},
	'{9,0,0,0,9}

};
	
	
	
	five <= '{

	'{9,9,9,9,9},
	'{9,0,0,0,0},
	'{9,9,9,9,9},
	'{0,0,0,0,9},
	'{9,9,9,9,9}

	};
	
	
	
	
	six <= '{
	
	'{9,9,9,9,9},
	'{9,0,0,0,9},
	'{9,9,9,9,9},
	'{0,0,0,0,9},
	'{9,9,9,9,9}

};
	
	
	
	
	seven <= '{
	
	'{9,0,0,0,0},
	'{9,0,0,0,0},
	'{9,0,0,0,0},
	'{9,0,0,0,9},
	'{9,9,9,9,9}

};

	eight <= '{
	
	'{9,9,9,9,9},
	'{9,0,0,0,9},
	'{9,9,9,9,9},
	'{9,0,0,0,9},
	'{9,9,9,9,9}


};	
	
	nine <= '{
	
	'{9,9,9,9,9},
	'{9,0,0,0,0},
	'{9,9,9,9,9},
	'{9,0,0,0,9},
	'{9,9,9,9,9}

};
	
ANNWU <= '{

		'{9,9,9,9,9,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,9,0,0,0,9,0,9,0,0,0,9},
		'{9,0,0,0,9,0,9,9,0,9,9,0,0,0,9,9,0,0,9,0,9,9,0,0,9,0,9,0,0,0,9},
		'{9,0,0,0,9,0,9,0,9,0,9,0,0,0,9,0,9,0,9,0,9,0,9,0,9,0,9,9,9,9,9},
		'{9,0,0,0,9,0,9,0,0,0,9,0,0,0,9,0,0,9,9,0,9,0,0,9,9,0,9,0,0,0,9},
		'{9,0,0,0,9,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,9,0,0,0,9,0,9,9,9,9,9}
};

PATRICKSU <= '{

		'{9,9,9,9,9,0,9,9,9,9,9,0,0,0,9,0,0,9,0,9,9,9,9,9,0,9,9,9,9,9,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,0,0,0,0,9},
		'{9,0,0,0,9,0,9,0,0,0,0,0,0,0,0,9,0,9,0,0,0,0,0,9,0,0,0,9,0,0,0,0,9,0,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,0,0,0,0,9},
		'{9,0,0,0,9,0,9,9,9,9,9,0,0,0,0,0,9,9,0,0,0,0,0,9,0,0,0,9,0,0,0,9,9,9,9,9,0,0,0,9,0,0,0,9,9,9,9,9,0,9,9,9,9,9},
		'{9,0,0,0,9,0,0,0,0,0,9,0,0,0,0,9,0,9,0,0,0,0,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,0,0,9,0,9,0,0,0,9},
		'{9,0,0,0,9,0,9,9,9,9,9,0,0,0,9,0,0,9,0,9,9,9,9,9,0,9,9,9,9,9,0,9,9,9,9,9,0,9,9,9,9,9,0,9,9,9,9,9,0,9,9,9,9,9}
};
	end
endmodule 
	

