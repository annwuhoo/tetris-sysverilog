//Block Hard Way

module Sprite_Table (
					// variable [#Rows][#Cols][EntryDepth]
					 output logic [15:0][63:0][2:0] I_block_h,
					 output logic [63:0][15:0][2:0] I_block_v,
					 output logic [31:0][31:0][2:0] O_block);
					 // output logic [15:0][23:0][4:0] J_block_1,
//					 output logic [319:0][159:0][4:0] Board);
	
	//Single Standard Block is 16x16
	always_comb
	begin
//	 I_block_h <= '{
//		
//		//64 long and 16 high
//		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
//		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
//		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
//		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}
//
//		};


	 I_block_h <= '{
		
		//64 long and 16 high
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,2,2,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,2,2,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,2,2,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,2,2,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,2,2,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,2,2,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7,1,1,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}

		};
	
	I_block_v <= '{
	
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}, // 16 long
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}, // 64 high
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,1,1,1,1,1,1,1,1,1,1,1,1,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}
		
		};
	
	O_block <= '{
	
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}, // 32 long
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}, // 32 high
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
	   '{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
	   '{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
	   '{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
	   '{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
	   '{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
	   '{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
	   '{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
	   '{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7,7,7,2,2,2,2,2,2,2,2,2,2,2,2,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7},
		'{7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7,7}
	
	};
	
//	J_block_1 <= '{
//	
//		'{9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9}, //24 wide
//		'{9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9}, //16 high
//		'{9,3,3,3,3,3,3,9,9,3,3,3,3,3,9,9,3,3,3,3,3,3,3,9},
//		'{9,3,3,3,3,3,3,9,9,3,3,3,3,3,9,9,3,3,3,3,3,3,3,9},
//		'{9,3,3,3,3,3,3,9,9,3,3,3,3,3,9,9,3,3,3,3,3,3,3,9},
//		'{9,3,3,3,3,3,3,9,9,3,3,3,3,3,9,9,3,3,3,3,3,3,3,9},
//		'{9,3,3,3,3,3,3,9,9,3,3,3,3,3,9,9,3,3,3,3,3,3,3,9},
//		'{9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9},
//		'{9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9,9},
//		'{9,3,3,3,3,3,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
//		'{9,3,3,3,3,3,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
//		'{9,3,3,3,3,3,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
//		'{9,3,3,3,3,3,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
//		'{9,3,3,3,3,3,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
//		'{9,9,9,9,9,9,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0},
//		'{9,9,9,9,9,9,9,9,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0}
//
//		
//	};
	

	end
endmodule 